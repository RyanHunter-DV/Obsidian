`ifndef RhDebugger__sv
`define RhDebugger__sv
package RhDebugger;

	`include "uvm_macros.svh"
	import uvm_pkg::*;

	`include "rhlib.svh"
	`include "RhdMacros.svh"

	`include "RhdUserInterface.svh"

	// Log features
	`include "RhdInfoProcessor.svh"
	// TODO, no necessary, `include "RhdInfo.svh"
	// Thread features
	`include "threads/RhdThread.svh"
	`include "threads/RhdThreadProcessor.svh"
	// Breakpoint features
	`include "breakpoints/RhdBreakpoint.svh"
	`include "breakpoints/RhdBreakpointProcessor.svh"

	`include "RhdCore.svh"

endpackage


`endif



